//Aquí se realizará el auto chequeo de test bench